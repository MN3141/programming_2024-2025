library ieee;
use ieee.std_logic_1164.all; --include arrays

entity ent is

end ent;

architecture arch of ent is

begin

end arch;